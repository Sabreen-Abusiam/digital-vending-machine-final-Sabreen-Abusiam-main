// week5_ex2_mux_structural.v - 2-to-1 Multiplexer (Structural)
module week5_ex2_mux_structural(
 
);


endmodule
