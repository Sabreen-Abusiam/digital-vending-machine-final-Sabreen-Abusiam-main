// ex09.v - Overflow detection in addition
// WHAT TO DO: Detect when adding two numbers produces a result too large to fit in 5 bits.
// Overflow detection prevents errors when accumulating coins in the vending machine.
module ex09(
 
);


endmodule

