// ex12.v - POS form for payment check
// WHAT TO DO: Express the same logic function as Product of Sums (AND of ORs).
// You'll see that the same function can be written in different but equivalent ways.
module ex12(

);
 endmodule
