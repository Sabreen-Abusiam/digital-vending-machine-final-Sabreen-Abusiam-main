// ex14.v - Boolean theorems (De Morgan's, Absorption)
// WHAT TO DO: Apply De Morgan's theorem to convert between AND/OR operations with NOT.
// This powerful theorem lets you transform logic expressions to find simpler implementations.
module ex14(

);

 

endmodule

