// ex30.v - FSM state encoding (binary vs one-hot)
// WHAT TO DO: Learn two different ways to encode states - binary (fewer bits) and one-hot (faster).
// This shows you design tradeoffs between circuit size and speed.
module ex30(
  
);


endmodule

