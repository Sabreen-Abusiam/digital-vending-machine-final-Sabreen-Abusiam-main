// ex00.v - Your First Empty Verilog Moduleaa
// This verifies that your Verilog environment is set up correctly

module ex00();

  // This is an empty module - it does nothing!
  // But it's important to check that it compiles without errors
  
  // In real projects, you'll add inputs, outputs, and logic here
  // For now, this just tests that your Verilog tools work
  
endmodule
