// week5_ex3_truth_table_assign.v - Truth Table Implementation (Behavioral Assign)
module week5_ex3_truth_table_assign(
 
);


endmodule
