// ex10.v - Comparison circuit (paid >= price)
// WHAT TO DO: Build a comparator that checks if the customer paid enough for their product.
// This circuit outputs true when paid amount is greater than or equal to the price.
module ex10(
 
);



endmodule

