// ex47.v - RAM with read/write control
// WHAT TO DO: Add separate read and write enable signals for better memory control.
// This prevents accidental reads or writes by requiring explicit enable signals.
module ex47(

);


endmodule

