// week5_ex1_xor_always.v - XOR Gate (Behavioral Always)
module week5_ex1_xor_always(
 
);


endmodule
