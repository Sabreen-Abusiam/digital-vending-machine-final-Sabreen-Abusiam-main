// ex48.v - ROM for product prices
// WHAT TO DO: Create Read-Only Memory that stores fixed product prices.
// ROM is perfect for constant data that never changes, like price lists.
module ex48(
  
);



endmodule

