// week5_ex1_or_assign.v - OR Gate (Behavioral Assign)
module week5_ex1_or_assign(
 
);


endmodule
