// week5_ex6_challenge_circuit_assign.v - Challenge Circuit (Behavioral Assign)
module week5_ex6_challenge_circuit_assign(
 
);


endmodule
