// week5_ex1_not_assign.v - NOT Gate (Behavioral Assign)
module week5_ex1_not_assign(
 
);


endmodule
