// week5_ex1_nand_assign.v - NAND Gate (Behavioral Assign)
module week5_ex1_nand_assign(
 
);


endmodule
