// week5_ex1_nor_assign.v - NOR Gate (Behavioral Assign)
module week5_ex1_nor_assign(
 
);


endmodule
