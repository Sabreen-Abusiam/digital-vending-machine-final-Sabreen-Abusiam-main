// week5_ex2_encoder_always.v - 4-to-2 Encoder (Behavioral Always)
module week5_ex2_encoder_always(
 
);


endmodule
