// week5_ex4_simple_circuit_assign.v - Simple Circuit (Behavioral Assign)
module week5_ex4_simple_circuit_assign(
 
);


endmodule
