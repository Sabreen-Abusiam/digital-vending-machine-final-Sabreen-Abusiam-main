// ex06.v - Binary Addition (Adding Two Coins)
// This demonstrates multi-bit signals and arithmetic operations

module ex06(
  
endmodule
