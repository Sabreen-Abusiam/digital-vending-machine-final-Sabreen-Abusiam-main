// ex11.v - SOP form for payment check
// WHAT TO DO: Express a logic function as Sum of Products (OR of ANDs).
// This teaches you one standard way to write Boolean expressions used in digital design.
module ex11(

);

  // F = A'B'C + A'BC = A'C(B' + B) = A'C
 

endmodule

