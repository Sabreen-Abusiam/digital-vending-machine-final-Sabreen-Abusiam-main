// week5_ex1_nand_always.v - NAND Gate (Behavioral Always)
module week5_ex1_nand_always(
 
);


endmodule
