// ex46.v - Simple RAM (4 locations, 4-bit data)
// WHAT TO DO: Create your first Random Access Memory to store and retrieve data.
// RAM uses an address to select which location to read from or write to.
module ex46(
 
);

9

endmodule

