// ex50.v - Complete Vending Machine System (Final Integration)
// WHAT TO DO: Integrate ALL concepts into one complete working vending machine!
// This is your final project combining FSM, arithmetic, memory, and all skills you've learned.

// ALU module for arithmetic operations
module alu_vending(

);


endmodule

