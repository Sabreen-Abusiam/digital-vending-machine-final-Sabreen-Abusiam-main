// ex43.v - ALU with comparison (CMP)
// WHAT TO DO: Add comparison operations that output flags for equal and greater-than.
// These flags are used for decision making in the vending machine controller.
module ex43(

);


endmodule

