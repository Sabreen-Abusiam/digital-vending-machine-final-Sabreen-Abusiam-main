// week5_ex5_advanced_circuit_structural.v - Advanced Circuit (Structural)
module week5_ex5_advanced_circuit_structural(
 
);


endmodule
