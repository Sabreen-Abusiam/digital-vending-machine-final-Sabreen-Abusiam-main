// ex26.v - Simple 2-State Finite State Machine (FSM)
// FSMs are used to control sequences of operations
// Like a traffic light or vending machine controller

module ex26(

);

  // States: 0 = IDLE, 1 = ACTIVE

endmodule
