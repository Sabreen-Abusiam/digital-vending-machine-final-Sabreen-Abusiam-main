// ex49.v - Inventory management with RAM
// WHAT TO DO: Use RAM to track product inventory, decrementing stock when items are dispensed.
// This adds realistic inventory management to your vending machine.
module ex49(
  
);

endmodule

