// ex27.v - 3-state FSM (IDLE, ACCEPT, CHECK)
// WHAT TO DO: Expand your FSM to three states to handle coin acceptance and checking.
// This teaches you how FSMs transition through multiple states based on inputs.
module ex27(

);


endmodule

