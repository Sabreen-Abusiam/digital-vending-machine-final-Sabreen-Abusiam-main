// week5_ex3_truth_table_structural.v - Truth Table Implementation (Structural)
module week5_ex3_truth_table_structural(
 
);


endmodule
