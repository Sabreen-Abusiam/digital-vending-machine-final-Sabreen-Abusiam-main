// week5_ex1_and_assign.v - AND Gate (Behavioral Assign)
module week5_ex1_and_assign(
 
);


endmodule
