// week5_ex2_encoder_assign.v - 4-to-2 Encoder (Behavioral Assign)
module week5_ex2_encoder_assign(
 
);


endmodule
