// week5_ex2_encoder_structural.v - 4-to-2 Encoder (Structural)
module week5_ex2_encoder_structural(
 
);


endmodule

