// ex38.v - 4-bit ripple-carry adder
// WHAT TO DO: Chain multiple full adders together to create a 4-bit adder circuit.
// Ripple-carry means the carry "ripples" from bit 0 to bit 3 sequentially.
module ex38(

);



endmodule

