// week5_ex1_or_always.v - OR Gate (Behavioral Always)
module week5_ex1_or_always(
 
);


endmodule
