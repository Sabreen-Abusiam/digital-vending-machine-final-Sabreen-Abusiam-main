// week5_ex3_truth_table_always.v - Truth Table Implementation (Behavioral Always)
module week5_ex3_truth_table_always(
 
);


endmodule
