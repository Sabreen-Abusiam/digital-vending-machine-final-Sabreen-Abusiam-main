// ex15.v - Consensus theorem
// WHAT TO DO: Use the consensus theorem to eliminate redundant terms in Boolean expressions.
// This optimization reduces the number of gates needed in your circuit.
module ex15(
 
);


endmodule

