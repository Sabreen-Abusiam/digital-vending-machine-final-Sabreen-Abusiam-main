// ex19.v - 2:1 and 4:1 Multiplexers
// WHAT TO DO: Build a multiplexer (MUX) that selects one input from multiple options.
// MUXes are like digital switches - select signals choose which input passes to output.
module ex19(

);

  // 4:1 MUX: Y = D[sel]


endmodule

