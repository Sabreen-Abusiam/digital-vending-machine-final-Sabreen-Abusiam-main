// week5_ex2_mux_always.v - 2-to-1 Multiplexer (Behavioral Always)
module week5_ex2_mux_always(
 
);


endmodule
