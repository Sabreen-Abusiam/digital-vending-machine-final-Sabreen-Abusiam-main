// ex33.v - Product dispenser FSM
// WHAT TO DO: Build a controlled dispenser that only releases products when payment is confirmed.
// This prevents giving away free products - dispense only when both request AND payment are valid.
module ex33(

);



endmodule

