// week5_ex1_xor_assign.v - XOR Gate (Behavioral Assign)
module week5_ex1_xor_assign(
 
);


endmodule
