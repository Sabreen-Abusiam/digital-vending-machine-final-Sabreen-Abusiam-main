// week5_ex2_decoder_structural.v - 2-to-4 Decoder (Structural)
module week5_ex2_decoder_structural(
 
);


endmodule
