// ex31.v - Coin accumulator with FSM
// WHAT TO DO: Combine sequential logic (register) with FSM to accumulate coin values.
// This integrates your register from Part 5 with state machine control to track total money.
module ex31(

);

endmodule

