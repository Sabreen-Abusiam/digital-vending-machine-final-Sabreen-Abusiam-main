// week5_ex2_decoder_always.v - 2-to-4 Decoder (Behavioral Always)
module week5_ex2_decoder_always(
 
);


endmodule
