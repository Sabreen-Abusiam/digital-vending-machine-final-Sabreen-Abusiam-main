// ex34.v - Change calculator FSM
// WHAT TO DO: Implement a sequential circuit that calculates and stores the change to return.
// This uses a register to hold the change value (paid - price) until it's dispensed.
module ex34(

);

endmodule

