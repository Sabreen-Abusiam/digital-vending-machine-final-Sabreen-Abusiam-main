// ex35.v - Combinational logic using always @(*)
// WHAT TO DO: Learn to use always @(*) blocks for combinational logic with case statements.
// This is an alternative to assign statements, useful for complex multi-operation circuits.
module ex35(

);



endmodule

