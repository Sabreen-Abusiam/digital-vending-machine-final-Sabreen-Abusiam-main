// ex41.v - Simple 2-operation ALU (ADD/SUB)
// WHAT TO DO: Build your first Arithmetic Logic Unit that performs ADD or SUB based on opcode.
// ALUs are the computational heart of processors - this is a simplified version.
module ex41(
 
);



endmodule

