// ex40.v - Combined Adder/Subtractor unit
// WHAT TO DO: Create one circuit that can both add and subtract based on a control signal.
// This is more efficient than having separate adder and subtractor circuits.
module ex40(

);


endmodule

