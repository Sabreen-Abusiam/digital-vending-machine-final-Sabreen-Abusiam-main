// week5_ex6_challenge_circuit_structural.v - Challenge Circuit (Structural)
module week5_ex6_challenge_circuit_structural(
 
);


endmodule
