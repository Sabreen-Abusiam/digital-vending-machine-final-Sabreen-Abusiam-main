// week5_ex4_simple_circuit_structural.v - Simple Circuit (Structural)
module week5_ex4_simple_circuit_structural(
 
);


endmodule
