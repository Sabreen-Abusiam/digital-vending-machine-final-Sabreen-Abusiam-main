// week5_ex1_nor_always.v - NOR Gate (Behavioral Always)
module week5_ex1_nor_always(
 
);


endmodule
