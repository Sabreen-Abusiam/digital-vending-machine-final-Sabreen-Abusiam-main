// ex38.v - 4-bit ripple-carry adder
// WHAT TO DO: Chain multiple full adders together to create a 4-bit adder circuit.
// Ripple-carry means the carry "ripples" from bit 0 to bit 3 sequentially.
module ex38(
    input  [3:0] a,
    input  [3:0] b,
    input        cin,
    output [3:0] sum,
    output       cout
);

    wire c1, c2, c3;

    ex37 fa0(.a(a[0]), .b(b[0]), .cin(cin), .sum(sum[0]), .cout(c1));
    ex37 fa1(.a(a[1]), .b(b[1]), .cin(c1),  .sum(sum[1]), .cout(c2));
    ex37 fa2(.a(a[2]), .b(b[2]), .cin(c2),  .sum(sum[2]), .cout(c3));
    ex37 fa3(.a(a[3]), .b(b[3]), .cin(c3),  .sum(sum[3]), .cout(cout));

endmodule