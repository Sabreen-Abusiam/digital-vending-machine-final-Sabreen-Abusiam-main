// ex44.v - ALU with flags (carry, zero, negative)
// WHAT TO DO: Generate status flags that indicate properties of the ALU result.
// Carry (overflow), zero, and negative flags help detect special conditions.
module ex44(

);


endmodule

