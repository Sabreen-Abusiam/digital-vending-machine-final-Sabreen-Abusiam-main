// ex28.v - 4-state FSM for vending machine
// WHAT TO DO: Add a DISPENSE state to create a basic functioning vending machine controller.
// Now your FSM can accept coins, check payment, and dispense products.
module ex28(
 
);



endmodule


