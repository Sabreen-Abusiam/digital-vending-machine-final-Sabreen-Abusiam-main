// week5_ex1_and_always.v - AND Gate (Behavioral Always)
module week5_ex1_and_always(
 
);


endmodule
