// week5_soda_machine_fsm.v - Soda Machine FSM Controller
// Exercise 3.26: Design an FSM controller for a soda machine
// Sodas cost 25 cents. Machine accepts nickels (5¢), dimes (10¢), and quarters (25¢)
// When enough coins are inserted, dispenses soda and returns change
// Then ready to accept coins for another soda

module week5_soda_machine_fsm(
  
);


endmodule



