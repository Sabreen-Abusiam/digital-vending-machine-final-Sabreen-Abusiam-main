// week5_ex4_simple_circuit_always.v - Simple Circuit (Behavioral Always)
module week5_ex4_simple_circuit_always(
 
);


endmodule
