// ex29.v - 5-state complete FSM
// WHAT TO DO: Add a CHANGE state to complete the full vending machine transaction cycle.
// This final state handles returning change before going back to IDLE for the next customer.
module ex29(

);


endmodule

