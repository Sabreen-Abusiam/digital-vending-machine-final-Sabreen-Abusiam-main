// week5_ex6_challenge_circuit_always.v - Challenge Circuit (Behavioral Always)
module week5_ex6_challenge_circuit_always(
 
);


endmodule
