// week5_ex5_advanced_circuit_assign.v - Advanced Circuit (Behavioral Assign)
module week5_ex5_advanced_circuit_assign(
 
);


endmodule
