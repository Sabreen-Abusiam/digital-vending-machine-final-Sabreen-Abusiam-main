// ex42.v - 4-operation ALU (ADD/SUB/AND/OR)
// WHAT TO DO: Expand your ALU to perform four operations: arithmetic (ADD/SUB) and logic (AND/OR).
// Use a 2-bit opcode to select which operation to perform.
module ex42(

);


endmodule

