// ex39.v - 5-bit subtractor for change
// WHAT TO DO: Build a subtractor circuit to calculate change (paid - price).
// Subtraction can be implemented using addition with 2's complement.
module ex39(
 
);



endmodule

