// week5_ex2_mux_assign.v - 2-to-1 Multiplexer (Behavioral Assign)
module week5_ex2_mux_assign(
 
);


endmodule
