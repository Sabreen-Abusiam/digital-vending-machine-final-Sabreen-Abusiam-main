// ex32.v - Payment validator FSM
// WHAT TO DO: Create a clocked circuit that continuously checks if payment is sufficient.
// This validates that the customer has inserted enough money before allowing a purchase.
module ex32(

);


endmodule

