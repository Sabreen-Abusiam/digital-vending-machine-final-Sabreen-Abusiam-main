// ex45.v - Complete ALU with all operations
// WHAT TO DO: Build a full-featured ALU with 8 operations including shifts and XOR.
// This is similar to what you'd find in a real processor's arithmetic unit.
module ex45(

);



endmodule

