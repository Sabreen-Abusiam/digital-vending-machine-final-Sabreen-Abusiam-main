// week5_ex1_not_always.v - NOT Gate (Behavioral Always)
module week5_ex1_not_always(
 
);


endmodule
