// week5_ex2_decoder_assign.v - 2-to-4 Decoder (Behavioral Assign)
module week5_ex2_decoder_assign(
 
);


endmodule
