// week5_ex5_advanced_circuit_always.v - Advanced Circuit (Behavioral Always)
module week5_ex5_advanced_circuit_always(
 
);


endmodule
