// ex25.v - Register with load and clear
// WHAT TO DO: Combine load (enable) and clear (reset) controls in one register.
// This gives you full control over when to store new values and when to reset to zero.
module ex25(
 
);



endmodule

