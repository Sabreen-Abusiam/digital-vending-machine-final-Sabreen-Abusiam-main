// ex13.v - Boolean axioms (Identity, Null, Idempotent)
// WHAT TO DO: Learn the basic rules of Boolean algebra (A OR 0 = A, A AND 1 = A, etc.).
// These fundamental laws help you simplify complex logic circuits.
module ex13(

);


endmodule

